----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    17:42:44 01/08/2008
-- Design Name:
-- Module Name:    memory_int - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.std_logic_textio.all;
use std.textio.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memory_int is
   port ( clk  : in  std_logic;
          addr : in  std_logic_vector (10 downto 0);
          inp  : in  std_logic_vector (15 downto 0);
          outp : out std_logic_vector (15 downto 0);
          we   : in  std_logic);
end memory_int;


architecture Simulation of memory_int is
   type saveArray is array (0 to (2**addr'length-1)) of std_logic_vector(15 downto 0);
   signal data : saveArray := (others => (others => '0'));
begin

   mem_ctrl: process(clk)
      variable init : integer := 0;
      file inputfile : text open read_mode is "../memory.txt";
      variable inputline : line;
      variable inputval  : std_logic_vector(15 downto 0);
      variable address   : integer := 0;

   begin
      if init = 0 then
         while not endfile(inputfile) loop
            readline(inputfile, inputline);
            hread(inputline, inputval);
            data(address) <= inputval;
            address := address+1;
         end loop;
         init := 1;
      elsif rising_edge(clk) then
         if we = '1' then
            data(conv_integer(unsigned(addr))) <= inp;
            outp <= inp;
         else
            outp <= data(conv_integer(unsigned(addr)));
         end if;
      end if;
   end process mem_ctrl;
end Simulation;


architecture Synthesis of memory_int is
   type saveArray is array (0 to (2**addr'length-1)) of std_logic_vector(15 downto 0);
   signal data : saveArray := ( X"c008",
  X"c222",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"8230",
  X"b000",
  X"8231",
  X"b005",
  X"8282",
  X"b001",
  X"8229",
  X"9274",
  X"8227",
  X"9271",
  X"9272",
  X"9273",
  X"9274",
  X"9275",
  X"9276",
  X"9277",
  X"9278",
  X"9279",
  X"927a",
  X"927b",
  X"f159",
  X"8271",
  X"d01d",
  X"f023",
  X"8227",
  X"9271",
  X"c01d",
  X"8274",
  X"d041",
  X"8271",
  X"2234",
  X"d04c",
  X"8271",
  X"2235",
  X"d04f",
  X"8271",
  X"2236",
  X"d058",
  X"8271",
  X"2243",
  X"d05b",
  X"8271",
  X"2238",
  X"d07e",
  X"8271",
  X"2244",
  X"d095",
  X"8274",
  X"2228",
  X"d04b",
  X"8271",
  X"2239",
  X"e04b",
  X"8242",
  X"2271",
  X"e04b",
  X"c084",
  X"8271",
  X"2237",
  X"d06b",
  X"8271",
  X"2239",
  X"e04b",
  X"8242",
  X"2271",
  X"e04b",
  X"c084",
  X"a100",
  X"8227",
  X"9272",
  X"c052",
  X"8228",
  X"9272",
  X"c052",
  X"8227",
  X"9274",
  X"f0cc",
  X"8272",
  X"9278",
  X"c0a7",
  X"8228",
  X"9273",
  X"c05d",
  X"8229",
  X"9273",
  X"8227",
  X"9274",
  X"8279",
  X"d064",
  X"f0c1",
  X"827e",
  X"c065",
  X"8275",
  X"9277",
  X"8227",
  X"9275",
  X"8273",
  X"9279",
  X"c0a7",
  X"8227",
  X"9274",
  X"8276",
  X"b021",
  X"8277",
  X"b021",
  X"8278",
  X"b021",
  X"8279",
  X"b021",
  X"8227",
  X"9276",
  X"9277",
  X"9278",
  X"9279",
  X"827a",
  X"1228",
  X"927a",
  X"c0a7",
  X"827a",
  X"d04b",
  X"8228",
  X"9274",
  X"f0e4",
  X"c0a7",
  X"8229",
  X"9274",
  X"8275",
  X"927c",
  X"822a",
  X"927d",
  X"f0f3",
  X"8271",
  X"2239",
  X"127e",
  X"9275",
  X"a004",
  X"3232",
  X"d0a7",
  X"8228",
  X"927b",
  X"c0a7",
  X"827a",
  X"d099",
  X"f0e4",
  X"c095",
  X"f0cc",
  X"8276",
  X"9275",
  X"827b",
  X"d09f",
  X"c0a7",
  X"f184",
  X"8255",
  X"b002",
  X"f1b5",
  X"f1d3",
  X"f184",
  X"f1c8",
  X"c0af",
  X"827b",
  X"d0bd",
  X"f184",
  X"824f",
  X"b002",
  X"f1b5",
  X"f184",
  X"f1c8",
  X"8227",
  X"9275",
  X"9276",
  X"9277",
  X"9278",
  X"9279",
  X"927a",
  X"927b",
  X"9274",
  X"8229",
  X"9274",
  X"8282",
  X"b001",
  X"a100",
  X"8271",
  X"9281",
  X"f194",
  X"a100",
  X"8275",
  X"927d",
  X"8277",
  X"927c",
  X"8279",
  X"2228",
  X"d0ca",
  X"f11f",
  X"c0cb",
  X"f0f3",
  X"a100",
  X"8279",
  X"d0d3",
  X"f0c1",
  X"827e",
  X"9275",
  X"8227",
  X"9279",
  X"8278",
  X"d0d9",
  X"8276",
  X"2275",
  X"9276",
  X"c0dc",
  X"8276",
  X"1275",
  X"9276",
  X"a004",
  X"3232",
  X"d0e1",
  X"8228",
  X"927b",
  X"8227",
  X"9275",
  X"a100",
  X"f0cc",
  X"8276",
  X"9275",
  X"a031",
  X"9279",
  X"a031",
  X"9278",
  X"a031",
  X"9277",
  X"a031",
  X"9276",
  X"827a",
  X"2228",
  X"927a",
  X"a100",
  X"8227",
  X"927e",
  X"927f",
  X"827c",
  X"e0f9",
  X"c0fe",
  X"5000",
  X"927c",
  X"827f",
  X"4000",
  X"927f",
  X"827d",
  X"e101",
  X"c106",
  X"5000",
  X"927d",
  X"827f",
  X"4000",
  X"927f",
  X"827d",
  X"d116",
  X"3228",
  X"d10e",
  X"827c",
  X"127e",
  X"e11c",
  X"927e",
  X"827c",
  X"127c",
  X"927c",
  X"e11c",
  X"827d",
  X"7000",
  X"927d",
  X"c107",
  X"827f",
  X"d11b",
  X"827e",
  X"5000",
  X"927e",
  X"a100",
  X"8228",
  X"927b",
  X"a100",
  X"8227",
  X"927e",
  X"927f",
  X"827c",
  X"e125",
  X"c12a",
  X"5000",
  X"927c",
  X"827f",
  X"4000",
  X"927f",
  X"827d",
  X"e12d",
  X"c132",
  X"5000",
  X"927d",
  X"827f",
  X"4000",
  X"927f",
  X"8228",
  X"9280",
  X"827c",
  X"227d",
  X"e13e",
  X"827d",
  X"127d",
  X"927d",
  X"8280",
  X"1280",
  X"9280",
  X"c134",
  X"827d",
  X"7000",
  X"927d",
  X"8280",
  X"7000",
  X"9280",
  X"d153",
  X"827c",
  X"227d",
  X"e14c",
  X"927c",
  X"8280",
  X"127e",
  X"927e",
  X"827d",
  X"7000",
  X"927d",
  X"8280",
  X"7000",
  X"9280",
  X"c144",
  X"827f",
  X"d158",
  X"827e",
  X"5000",
  X"927e",
  X"a100",
  X"f171",
  X"f1c8",
  X"826b",
  X"b002",
  X"f1b5",
  X"f184",
  X"f1c8",
  X"f184",
  X"8239",
  X"9281",
  X"f194",
  X"823a",
  X"9281",
  X"f194",
  X"823b",
  X"9281",
  X"f194",
  X"823c",
  X"9281",
  X"f194",
  X"823d",
  X"9281",
  X"f194",
  X"a100",
  X"826c",
  X"b003",
  X"826d",
  X"9284",
  X"8246",
  X"b023",
  X"8284",
  X"2228",
  X"9284",
  X"d17c",
  X"c175",
  X"826c",
  X"9285",
  X"b003",
  X"8227",
  X"9286",
  X"8228",
  X"9287",
  X"a100",
  X"8228",
  X"9287",
  X"8227",
  X"9286",
  X"8285",
  X"126e",
  X"9285",
  X"b003",
  X"826f",
  X"2285",
  X"e190",
  X"a100",
  X"826c",
  X"9285",
  X"b003",
  X"a100",
  X"8287",
  X"d1ac",
  X"8281",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"9288",
  X"3248",
  X"b013",
  X"8227",
  X"9287",
  X"1286",
  X"9286",
  X"8270",
  X"2286",
  X"e1aa",
  X"a100",
  X"f184",
  X"a100",
  X"8281",
  X"1288",
  X"b023",
  X"8228",
  X"9287",
  X"8228",
  X"1286",
  X"9286",
  X"a100",
  X"a012",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"d1c7",
  X"9281",
  X"f194",
  X"a022",
  X"324a",
  X"d1c7",
  X"9281",
  X"f194",
  X"c1b5",
  X"a100",
  X"826e",
  X"9284",
  X"8245",
  X"b023",
  X"8284",
  X"2228",
  X"9284",
  X"d1d1",
  X"c1ca",
  X"f184",
  X"a100",
  X"8227",
  X"9289",
  X"928a",
  X"928b",
  X"928c",
  X"928d",
  X"8275",
  X"e21b",
  X"8275",
  X"222c",
  X"9275",
  X"e1e3",
  X"8289",
  X"1228",
  X"9289",
  X"c1db",
  X"122c",
  X"222d",
  X"9275",
  X"e1ec",
  X"828a",
  X"1228",
  X"928a",
  X"8275",
  X"c1e4",
  X"122d",
  X"222e",
  X"9275",
  X"e1f5",
  X"828b",
  X"1228",
  X"928b",
  X"8275",
  X"c1ed",
  X"122e",
  X"222f",
  X"9275",
  X"e1fe",
  X"828c",
  X"1228",
  X"928c",
  X"8275",
  X"c1f6",
  X"122f",
  X"928d",
  X"8289",
  X"d20c",
  X"f217",
  X"828a",
  X"f217",
  X"828b",
  X"f217",
  X"828c",
  X"f217",
  X"828a",
  X"f217",
  X"a100",
  X"828a",
  X"d20f",
  X"c204",
  X"828b",
  X"d212",
  X"c206",
  X"828c",
  X"d215",
  X"c208",
  X"828d",
  X"c20a",
  X"1247",
  X"9281",
  X"f194",
  X"a100",
  X"5000",
  X"9275",
  X"8235",
  X"9281",
  X"f194",
  X"8275",
  X"c1db",
  X"b030",
  X"8fff",
  X"9271",
  X"a020",
  X"a200",
  X"0000",
  X"0001",
  X"0002",
  X"000a",
  X"ff00",
  X"2710",
  X"03e8",
  X"0064",
  X"000a",
  X"07ff",
  X"0102",
  X"0008",
  X"00ff",
  X"002b",
  X"002d",
  X"002a",
  X"0028",
  X"0029",
  X"0030",
  X"0031",
  X"0032",
  X"0033",
  X"0034",
  X"0035",
  X"0036",
  X"0037",
  X"0038",
  X"0039",
  X"002f",
  X"003d",
  X"2d2d",
  X"2020",
  X"0030",
  X"ff20",
  X"ff00",
  X"00ff",
  X"4572",
  X"726f",
  X"7221",
  X"0000",
  X"024b",
  X"5265",
  X"7375",
  X"6c74",
  X"3a20",
  X"0000",
  X"0250",
  X"5765",
  X"6c63",
  X"6f6d",
  X"6520",
  X"746f",
  X"2074",
  X"6865",
  X"2075",
  X"6c74",
  X"696d",
  X"6174",
  X"6520",
  X"4c4d",
  X"4520",
  X"6361",
  X"6c63",
  X"756c",
  X"6174",
  X"6f72",
  X"2120",
  X"0000",
  X"0256",
  X"0800",
  X"0640",
  X"0028",
  X"0e40",
  X"004f",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0283",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0001",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  others => X"0000" );
begin

   mem_ctrl: process(clk)
   begin
      if rising_edge(clk) then
         if we = '1' then
            data(conv_integer(unsigned(addr))) <= inp;
            outp <= inp;
         else
            outp <= data(conv_integer(unsigned(addr)));
         end if;
      end if;
   end process mem_ctrl;
end Synthesis;







