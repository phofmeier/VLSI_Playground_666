----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:23:38 06/11/2017 
-- Design Name: 
-- Module Name:    charecterRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_arith.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity characterRAM is
port (pixel_clk  : in std_logic;
		clk        : in STD_LOGIC;
		we         : in  STD_LOGIC;
		pixel_en   : in STD_LOGIC;
		pixel_left   : in STD_LOGIC;
		address_read : in std_logic_vector(11 downto 0);
		addressbus  : in std_logic_vector(11 downto 0);
		databus    : in  STD_LOGIC_VECTOR (15 downto 0);
		dataout    : out  STD_LOGIC_VECTOR (15 downto 0)); 
end characterRAM;	

architecture Behavioral of characterRAM is


type character_memory is array (0 to 1599) of std_logic_vector(15 downto 0);
 
signal VGA_RAM: character_memory:=
(X"2031",
X"5620",
X"534C",
X"2049",
X"6C50",
X"7961",
X"7267",
X"756F",
X"646E",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2032",
X"5620",
X"534C",
X"2049",
X"6C50",
X"7961",
X"7267",
X"756F",
X"646E",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2033",
X"5620",
X"534C",
X"2049",
X"6C50",
X"7961",
X"7267",
X"756F",
X"646E",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2061",
X"6161",
X"6161",
X"2020",
X"2020",
X"2061",
X"6161",
X"6120",
X"6161",
X"6161",
X"2020",
X"2020",
X"6161",
X"6161",
X"2061",
X"6161",
X"6120",
X"2020",
X"2020",
X"2020",
X"2061",
X"6161",
X"6161",
X"2020",
X"2e61",
X"6161",
X"6161",
X"2e20",
X"2020",
X"2020",
X"2e61",
X"2020",
X"2020",
X"2e61",
X"6161",
X"612e",
X"2020",
X"2020",
X"2020",
X"2020",
X"2060",
X"3838",
X"3827",
X"2020",
X"2020",
X"2060",
X"3838",
X"2720",
X"6038",
X"3838",
X"2020",
X"202e",
X"3850",
X"2720",
X"2060",
X"3838",
X"382e",
X"2020",
X"2020",
X"2020",
X"6438",
X"3838",
X"3827",
X"2038",
X"3838",
X"2720",
X"6059",
X"3838",
X"2e20",
X"6138",
X"3838",
X"2020",
X"2064",
X"3850",
X"2760",
X"5938",
X"6220",
X"2020",
X"2020",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"3838",
X"2020",
X"2038",
X"3838",
X"2020",
X"6438",
X"2720",
X"2020",
X"2020",
X"3838",
X"3838",
X"6220",
X"2020",
X"2064",
X"5027",
X"7c38",
X"3820",
X"2038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2038",
X"3838",
X"2020",
X"3838",
X"3820",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"3838",
X"2020",
X"2038",
X"3838",
X"3838",
X"5b20",
X"2020",
X"2020",
X"2020",
X"3838",
X"2059",
X"3838",
X"2e20",
X"6450",
X"2020",
X"7c38",
X"3820",
X"2020",
X"6056",
X"6261",
X"6164",
X"3838",
X"3820",
X"2038",
X"3838",
X"2020",
X"3838",
X"3820",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"3838",
X"2020",
X"2038",
X"3838",
X"6038",
X"3862",
X"2e20",
X"2020",
X"2020",
X"3838",
X"2020",
X"6038",
X"3838",
X"2720",
X"2020",
X"7c38",
X"3820",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2720",
X"2038",
X"3838",
X"2020",
X"3838",
X"3820",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"6038",
X"382e",
X"2020",
X"2020",
X"2064",
X"3827",
X"2020",
X"2038",
X"3838",
X"2020",
X"6038",
X"3862",
X"2e20",
X"2020",
X"3838",
X"2020",
X"2020",
X"5920",
X"2020",
X"2020",
X"7c38",
X"3820",
X"2020",
X"2020",
X"202e",
X"3838",
X"5027",
X"2020",
X"2038",
X"3838",
X"2020",
X"6038",
X"3862",
X"2020",
X"6438",
X"3827",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"6059",
X"6261",
X"6164",
X"5027",
X"2020",
X"2020",
X"6138",
X"3838",
X"6120",
X"2061",
X"3838",
X"3861",
X"2061",
X"3838",
X"6120",
X"2020",
X"2020",
X"2020",
X"2061",
X"3838",
X"3861",
X"2020",
X"202e",
X"6150",
X"2720",
X"2020",
X"2020",
X"6138",
X"3838",
X"6120",
X"2060",
X"5938",
X"6264",
X"3850",
X"2720",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"3d3d",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2e64",
X"3838",
X"3838",
X"3862",
X"2e20",
X"2020",
X"2020",
X"2020",
X"2020",
X"2064",
X"3838",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2020",
X"2e64",
X"3838",
X"3838",
X"3862",
X"2e20",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2064",
X"3838",
X"5020",
X"2020",
X"5938",
X"3862",
X"2020",
X"2020",
X"2020",
X"2020",
X"6438",
X"3838",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2064",
X"3838",
X"5020",
X"2020",
X"5938",
X"3862",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2064",
X"3838",
X"5038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"6438",
X"3850",
X"2038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2064",
X"3838",
X"5020",
X"2038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"6438",
X"3850",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3820",
X"2020",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2059",
X"3838",
X"6220",
X"2020",
X"6438",
X"3850",
X"2020",
X"2064",
X"3838",
X"3838",
X"3838",
X"3838",
X"3838",
X"2020",
X"2020",
X"3838",
X"3861",
X"6161",
X"6161",
X"2020",
X"2059",
X"3838",
X"6220",
X"2020",
X"6438",
X"3850",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2259",
X"3838",
X"3838",
X"3850",
X"2220",
X"2020",
X"6438",
X"3850",
X"2020",
X"2020",
X"2038",
X"3838",
X"2020",
X"2020",
X"3838",
X"3838",
X"3838",
X"3838",
X"2020",
X"2020",
X"2259",
X"3838",
X"3838",
X"3850",
X"2220",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020",
X"2020");

begin

process(databus,addressbus,we,clk)
begin
	if (rising_edge(clk)) then 
		if (we = '1') then 
			VGA_RAM(conv_integer(addressbus))<=databus;
		end if;
	end if;
end process;

process(address_read,pixel_en,pixel_clk)
begin	
		if((pixel_en='1')) then 
			dataout<= VGA_RAM(conv_integer(address_read));
		else
			dataout <="ZZZZZZZZZZZZZZZZ";
		end if;
end process;
														
end Behavioral;

