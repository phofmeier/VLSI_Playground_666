library ieee;
use ieee.std_logic_1164.all;

package fontROM is

  type fontROMArray is array (0 to 256*12-1) of std_logic_vector(7 downto 0);  -- array definition for font ROM

  constant fontROM : fontROMArray := ( X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"08", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"30", X"0c", X"00", X"03", X"1c", X"00", X"0c", X"00", X"03", X"00", X"08", X"06", X"00", X"1e", X"30", X"00", X"00", X"0c", X"00", X"03", X"0c", X"03", X"00", X"00", X"33", X"00", X"3c", X"00", X"00", X"70", X"30", X"30", X"30", X"30", X"00", X"6e", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"24", X"aa", X"b6", X"18", X"18", X"30", X"1e", X"06", X"00", X"66", X"66", X"00", X"66", X"00", X"33", X"00", X"18", X"18", X"00", X"18", X"00", X"18", X"00", X"6e", X"66", X"00", X"66", X"00", X"66", X"00", X"66", X"00", X"33", X"00", X"1e", X"00", X"06", X"00", X"18", X"1e", X"00", X"18", X"00", X"ff", X"00", X"00", X"06", X"ff", X"18", X"00", X"1e", X"06", X"00", X"6e", X"00", X"00", X"00", X"18", X"1e", X"06", X"60", X"18", X"00", X"30", X"00", X"00", X"00", X"07", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                                       X"00", X"7e", X"7e", X"00", X"08", X"18", X"18", X"00", X"00", X"00", X"00", X"7c", X"3c", X"00", X"fe", X"00", X"01", X"40", X"18", X"66", X"fe", X"7e", X"00", X"18", X"18", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"66", X"36", X"0c", X"00", X"0e", X"0c", X"30", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"3e", X"08", X"1e", X"1e", X"30", X"3f", X"1c", X"7f", X"1e", X"1e", X"00", X"00", X"30", X"00", X"06", X"1e", X"3e", X"0c", X"3f", X"3c", X"1f", X"7f", X"7f", X"3c", X"33", X"1e", X"78", X"67", X"0f", X"63", X"63", X"1c", X"3f", X"1c", X"3f", X"1e", X"3f", X"33", X"33", X"63", X"33", X"33", X"7f", X"3c", X"00", X"3c", X"1c", X"00", X"0c", X"00", X"07", X"00", X"38", X"00", X"1c", X"00", X"07", X"18", X"30", X"07", X"1e", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"38", X"18", X"07", X"ce", X"00", X"1e", X"33", X"18", X"1e", X"33", X"06", X"36", X"00", X"1e", X"33", X"06", X"36", X"1c", X"0c", X"33", X"33", X"18", X"00", X"7c", X"1e", X"33", X"06", X"1e", X"06", X"66", X"33", X"00", X"00", X"66", X"5c", X"00", X"e8", X"18", X"18", X"18", X"18", X"6e", X"3b", X"1e", X"1e", X"0c", X"1c", X"00", X"46", X"c6", X"0c", X"00", X"00", X"49", X"55", X"eb", X"18", X"18", X"18", X"33", X"0c", X"1c", X"66", X"66", X"00", X"66", X"0c", X"33", X"00", X"18", X"18", X"00", X"18", X"00", X"18", X"6e", X"3b", X"66", X"00", X"66", X"00", X"66", X"00", X"66", X"00", X"0c", X"1f", X"33", X"33", X"0c", X"0f", X"0c", X"33", X"33", X"18", X"00", X"ff", X"00", X"18", X"0c", X"ff", X"0c", X"1e", X"33", X"0c", X"6e", X"3b", X"00", X"00", X"0f", X"0c", X"33", X"0c", X"30", X"0c", X"3f", X"18", X"00", X"00", X"00", X"cc", X"fe", X"7e", X"00", X"00", X"3c", X"33", X"00", X"0c", X"1e", X"1e", X"00", X"00",
                                       X"00", X"c3", X"ff", X"22", X"1c", X"3c", X"3c", X"00", X"00", X"00", X"00", X"70", X"66", X"00", X"c6", X"18", X"03", X"60", X"3c", X"66", X"eb", X"c6", X"00", X"3c", X"3c", X"18", X"00", X"00", X"00", X"00", X"08", X"7f", X"00", X"1e", X"66", X"36", X"3e", X"00", X"1b", X"0c", X"18", X"0c", X"00", X"00", X"00", X"00", X"00", X"40", X"63", X"0c", X"33", X"33", X"38", X"03", X"06", X"63", X"33", X"33", X"00", X"00", X"18", X"00", X"0c", X"33", X"63", X"1e", X"66", X"66", X"36", X"46", X"66", X"66", X"33", X"0c", X"30", X"66", X"06", X"77", X"63", X"36", X"66", X"36", X"66", X"33", X"2e", X"33", X"33", X"63", X"33", X"33", X"73", X"0c", X"01", X"30", X"36", X"00", X"18", X"00", X"06", X"00", X"30", X"00", X"36", X"00", X"06", X"18", X"30", X"06", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"04", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"18", X"0c", X"5b", X"00", X"33", X"33", X"0c", X"33", X"33", X"0c", X"36", X"00", X"33", X"33", X"0c", X"36", X"36", X"18", X"00", X"33", X"00", X"00", X"1e", X"33", X"33", X"0c", X"33", X"0c", X"66", X"00", X"33", X"00", X"06", X"36", X"00", X"18", X"0c", X"0c", X"0c", X"0c", X"3b", X"00", X"33", X"33", X"0c", X"22", X"00", X"67", X"67", X"0c", X"00", X"00", X"92", X"aa", X"6e", X"18", X"18", X"00", X"00", X"00", X"22", X"66", X"66", X"00", X"66", X"0c", X"33", X"00", X"18", X"18", X"00", X"18", X"00", X"18", X"3b", X"00", X"66", X"00", X"66", X"00", X"66", X"00", X"66", X"00", X"1b", X"36", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"18", X"00", X"ff", X"00", X"18", X"00", X"ff", X"00", X"33", X"00", X"00", X"3b", X"00", X"00", X"07", X"06", X"00", X"00", X"00", X"18", X"00", X"00", X"0c", X"00", X"0c", X"00", X"66", X"eb", X"c6", X"0c", X"00", X"66", X"00", X"00", X"0e", X"30", X"30", X"00", X"00",
                                       X"00", X"81", X"ff", X"77", X"3e", X"3c", X"7e", X"00", X"00", X"00", X"00", X"5c", X"66", X"00", X"fe", X"eb", X"07", X"70", X"7e", X"66", X"eb", X"0c", X"00", X"7e", X"7e", X"18", X"18", X"0c", X"00", X"24", X"08", X"7f", X"00", X"1e", X"66", X"7f", X"03", X"23", X"1b", X"0c", X"0c", X"18", X"66", X"18", X"00", X"00", X"00", X"60", X"73", X"0f", X"33", X"30", X"3c", X"03", X"03", X"63", X"33", X"33", X"1c", X"1c", X"0c", X"00", X"18", X"30", X"63", X"33", X"66", X"63", X"66", X"06", X"46", X"63", X"33", X"0c", X"30", X"36", X"06", X"7f", X"67", X"63", X"66", X"63", X"66", X"33", X"0c", X"33", X"33", X"63", X"33", X"33", X"19", X"0c", X"03", X"30", X"63", X"00", X"00", X"00", X"06", X"00", X"30", X"00", X"06", X"00", X"06", X"00", X"00", X"06", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"18", X"0c", X"73", X"08", X"33", X"00", X"00", X"00", X"00", X"00", X"1c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"1e", X"3f", X"00", X"1b", X"00", X"00", X"00", X"00", X"00", X"00", X"1e", X"33", X"00", X"06", X"73", X"00", X"18", X"00", X"00", X"00", X"00", X"00", X"63", X"33", X"33", X"00", X"5e", X"00", X"36", X"36", X"00", X"00", X"00", X"24", X"55", X"b6", X"18", X"18", X"0c", X"0c", X"0c", X"5e", X"66", X"66", X"00", X"66", X"1e", X"33", X"00", X"18", X"18", X"00", X"18", X"00", X"18", X"00", X"0c", X"66", X"00", X"66", X"00", X"66", X"00", X"66", X"00", X"30", X"66", X"3f", X"3f", X"3f", X"0c", X"1e", X"1e", X"1e", X"18", X"00", X"ff", X"00", X"18", X"1e", X"ff", X"1e", X"33", X"1e", X"1e", X"00", X"1e", X"00", X"06", X"3e", X"33", X"33", X"33", X"00", X"33", X"00", X"00", X"00", X"0c", X"00", X"3c", X"eb", X"0c", X"0c", X"00", X"66", X"00", X"00", X"0c", X"1c", X"18", X"3f", X"00",
                                       X"00", X"a5", X"db", X"7f", X"7f", X"ff", X"ff", X"00", X"00", X"00", X"00", X"4e", X"66", X"00", X"c6", X"7e", X"1f", X"7c", X"18", X"66", X"eb", X"3c", X"00", X"18", X"18", X"18", X"30", X"06", X"03", X"66", X"1c", X"3e", X"00", X"1e", X"24", X"36", X"03", X"33", X"0e", X"06", X"06", X"30", X"3c", X"18", X"00", X"00", X"00", X"30", X"7b", X"0c", X"30", X"30", X"36", X"03", X"03", X"60", X"33", X"33", X"1c", X"1c", X"06", X"7e", X"30", X"18", X"7b", X"33", X"66", X"03", X"66", X"26", X"26", X"03", X"33", X"0c", X"30", X"36", X"06", X"7f", X"6f", X"63", X"66", X"63", X"66", X"03", X"0c", X"33", X"33", X"63", X"1e", X"33", X"18", X"0c", X"06", X"30", X"00", X"00", X"00", X"1e", X"3e", X"1e", X"3e", X"1e", X"06", X"6e", X"36", X"1e", X"3c", X"66", X"18", X"3f", X"1f", X"1e", X"3b", X"6e", X"37", X"1e", X"3f", X"33", X"33", X"63", X"63", X"66", X"3f", X"06", X"18", X"18", X"00", X"1c", X"03", X"33", X"1e", X"1e", X"1e", X"1e", X"1f", X"1e", X"1e", X"1e", X"1e", X"1e", X"1e", X"1e", X"1e", X"1e", X"23", X"7f", X"1b", X"1e", X"1e", X"1e", X"33", X"33", X"66", X"33", X"33", X"1e", X"06", X"6b", X"00", X"7e", X"1e", X"1e", X"1e", X"33", X"1f", X"67", X"7e", X"1e", X"0c", X"55", X"00", X"1e", X"1e", X"0c", X"cc", X"33", X"49", X"aa", X"eb", X"18", X"18", X"1e", X"1e", X"1e", X"45", X"67", X"66", X"7f", X"67", X"33", X"1e", X"00", X"18", X"18", X"00", X"18", X"00", X"18", X"1e", X"1e", X"e6", X"fe", X"e7", X"ff", X"e6", X"ff", X"e7", X"00", X"60", X"66", X"23", X"23", X"23", X"0c", X"0c", X"0c", X"0c", X"18", X"00", X"ff", X"00", X"18", X"0c", X"ff", X"33", X"1b", X"33", X"33", X"1e", X"33", X"66", X"3e", X"66", X"33", X"33", X"33", X"66", X"33", X"00", X"00", X"00", X"3f", X"00", X"1f", X"eb", X"3c", X"00", X"00", X"66", X"00", X"00", X"0c", X"30", X"0c", X"3f", X"00",
                                       X"00", X"81", X"ff", X"7f", X"7f", X"e7", X"ff", X"00", X"00", X"00", X"00", X"1f", X"3c", X"00", X"c6", X"e7", X"7f", X"7f", X"18", X"66", X"ee", X"66", X"00", X"18", X"18", X"18", X"7f", X"7f", X"03", X"ff", X"1c", X"3e", X"00", X"0c", X"00", X"36", X"1e", X"18", X"5f", X"00", X"06", X"30", X"ff", X"7e", X"00", X"7f", X"00", X"18", X"6b", X"0c", X"18", X"1c", X"33", X"1f", X"1f", X"30", X"1e", X"3e", X"00", X"00", X"03", X"00", X"60", X"0c", X"7b", X"33", X"3e", X"03", X"66", X"3e", X"3e", X"03", X"3f", X"0c", X"30", X"1e", X"06", X"6b", X"7f", X"63", X"3e", X"63", X"3e", X"0e", X"0c", X"33", X"33", X"6b", X"0c", X"1e", X"0c", X"0c", X"0c", X"30", X"00", X"00", X"00", X"30", X"66", X"33", X"33", X"33", X"1f", X"33", X"6e", X"18", X"30", X"36", X"18", X"6b", X"33", X"33", X"66", X"33", X"76", X"33", X"06", X"33", X"33", X"63", X"36", X"66", X"31", X"03", X"00", X"30", X"00", X"36", X"03", X"33", X"33", X"30", X"30", X"30", X"30", X"33", X"33", X"33", X"33", X"18", X"18", X"18", X"33", X"33", X"03", X"e8", X"7f", X"33", X"33", X"33", X"33", X"33", X"66", X"33", X"33", X"33", X"3f", X"6b", X"63", X"18", X"30", X"18", X"33", X"33", X"33", X"6f", X"00", X"00", X"06", X"5e", X"3f", X"0c", X"ec", X"0c", X"66", X"66", X"92", X"55", X"6e", X"18", X"1f", X"33", X"33", X"33", X"45", X"60", X"66", X"60", X"60", X"03", X"3f", X"1f", X"f8", X"ff", X"ff", X"f8", X"ff", X"ff", X"30", X"33", X"06", X"06", X"00", X"00", X"06", X"00", X"00", X"63", X"7e", X"6f", X"03", X"03", X"03", X"3f", X"0c", X"0c", X"0c", X"1f", X"f8", X"ff", X"00", X"00", X"0c", X"ff", X"33", X"33", X"33", X"33", X"33", X"33", X"66", X"66", X"66", X"33", X"33", X"33", X"66", X"33", X"00", X"00", X"3f", X"0c", X"1f", X"ec", X"ee", X"66", X"3f", X"00", X"3c", X"00", X"18", X"1e", X"1e", X"3e", X"3f", X"00",
                                       X"00", X"bd", X"c3", X"7f", X"3e", X"e7", X"7e", X"00", X"00", X"00", X"00", X"33", X"18", X"00", X"c6", X"e7", X"1f", X"7c", X"18", X"00", X"e8", X"66", X"00", X"18", X"18", X"18", X"30", X"06", X"03", X"66", X"3e", X"1c", X"00", X"0c", X"00", X"36", X"30", X"0c", X"7b", X"00", X"06", X"30", X"3c", X"18", X"00", X"00", X"00", X"0c", X"6f", X"0c", X"0c", X"30", X"7f", X"30", X"33", X"18", X"33", X"18", X"00", X"00", X"06", X"7e", X"30", X"0c", X"7b", X"3f", X"66", X"03", X"66", X"26", X"26", X"73", X"33", X"0c", X"33", X"36", X"46", X"63", X"7b", X"63", X"06", X"73", X"36", X"18", X"0c", X"33", X"33", X"6b", X"1e", X"0c", X"06", X"0c", X"18", X"30", X"00", X"00", X"00", X"3e", X"66", X"03", X"33", X"3f", X"06", X"33", X"66", X"18", X"30", X"1e", X"18", X"6b", X"33", X"33", X"66", X"33", X"6e", X"06", X"06", X"33", X"33", X"6b", X"1c", X"66", X"18", X"06", X"18", X"18", X"00", X"63", X"03", X"33", X"3f", X"3e", X"3e", X"3e", X"3e", X"03", X"3f", X"3f", X"3f", X"18", X"18", X"18", X"33", X"33", X"1f", X"fe", X"1b", X"33", X"33", X"33", X"33", X"33", X"66", X"33", X"33", X"3b", X"06", X"6b", X"36", X"18", X"3e", X"18", X"33", X"33", X"33", X"7b", X"7f", X"7f", X"03", X"4e", X"30", X"76", X"f6", X"1e", X"33", X"cc", X"24", X"aa", X"b6", X"18", X"18", X"33", X"33", X"33", X"45", X"60", X"66", X"60", X"60", X"03", X"0c", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"3e", X"33", X"06", X"06", X"00", X"00", X"06", X"00", X"00", X"3e", X"63", X"66", X"1f", X"1f", X"1f", X"00", X"0c", X"0c", X"0c", X"00", X"18", X"ff", X"ff", X"18", X"0c", X"00", X"33", X"33", X"33", X"33", X"33", X"33", X"66", X"66", X"66", X"33", X"33", X"33", X"66", X"1e", X"00", X"00", X"00", X"0c", X"00", X"f6", X"e8", X"66", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3f", X"00",
                                       X"00", X"99", X"e7", X"3e", X"1c", X"18", X"18", X"00", X"00", X"00", X"00", X"33", X"7e", X"00", X"e6", X"7e", X"07", X"70", X"7e", X"00", X"e8", X"3c", X"7f", X"7e", X"18", X"7e", X"18", X"0c", X"7f", X"24", X"3e", X"1c", X"00", X"00", X"00", X"7f", X"30", X"06", X"33", X"00", X"0c", X"18", X"66", X"18", X"00", X"00", X"00", X"06", X"67", X"0c", X"06", X"30", X"30", X"30", X"33", X"0c", X"33", X"18", X"1c", X"1c", X"0c", X"00", X"18", X"00", X"03", X"33", X"66", X"63", X"66", X"06", X"06", X"63", X"33", X"0c", X"33", X"36", X"66", X"63", X"73", X"63", X"06", X"7b", X"66", X"33", X"0c", X"33", X"33", X"36", X"33", X"0c", X"46", X"0c", X"30", X"30", X"00", X"00", X"00", X"33", X"66", X"03", X"33", X"03", X"06", X"33", X"66", X"18", X"30", X"36", X"18", X"6b", X"33", X"33", X"66", X"33", X"06", X"18", X"06", X"33", X"33", X"6b", X"1c", X"66", X"06", X"0c", X"18", X"0c", X"00", X"63", X"33", X"33", X"03", X"33", X"33", X"33", X"33", X"03", X"03", X"03", X"03", X"18", X"18", X"18", X"3f", X"3f", X"03", X"1b", X"1b", X"33", X"33", X"33", X"33", X"33", X"66", X"33", X"33", X"37", X"06", X"67", X"1c", X"18", X"33", X"18", X"33", X"33", X"33", X"73", X"00", X"00", X"03", X"55", X"30", X"c3", X"eb", X"1e", X"33", X"cc", X"49", X"55", X"eb", X"18", X"18", X"3f", X"3f", X"3f", X"5e", X"67", X"66", X"67", X"7f", X"33", X"3f", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"33", X"3f", X"fe", X"e6", X"ff", X"e7", X"e6", X"ff", X"e7", X"36", X"63", X"66", X"03", X"03", X"03", X"00", X"0c", X"0c", X"0c", X"00", X"18", X"ff", X"ff", X"18", X"0c", X"00", X"33", X"33", X"33", X"33", X"33", X"33", X"66", X"3e", X"3e", X"33", X"33", X"33", X"66", X"0c", X"00", X"00", X"00", X"00", X"00", X"eb", X"e8", X"3c", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3f", X"00",
                                       X"00", X"c3", X"ff", X"1c", X"08", X"18", X"18", X"00", X"00", X"00", X"00", X"33", X"18", X"00", X"e7", X"eb", X"03", X"60", X"3c", X"66", X"e8", X"30", X"7f", X"3c", X"18", X"3c", X"00", X"00", X"00", X"00", X"7f", X"08", X"00", X"0c", X"00", X"36", X"1f", X"33", X"3b", X"00", X"18", X"0c", X"00", X"00", X"1c", X"00", X"1c", X"03", X"63", X"0c", X"33", X"33", X"30", X"33", X"33", X"0c", X"33", X"0c", X"1c", X"1c", X"18", X"00", X"0c", X"0c", X"03", X"33", X"66", X"66", X"36", X"46", X"06", X"66", X"33", X"0c", X"33", X"66", X"66", X"63", X"63", X"36", X"06", X"3e", X"66", X"33", X"0c", X"33", X"1e", X"36", X"33", X"0c", X"63", X"0c", X"60", X"30", X"00", X"00", X"00", X"33", X"66", X"33", X"33", X"33", X"06", X"3e", X"66", X"18", X"30", X"66", X"18", X"6b", X"33", X"33", X"66", X"33", X"06", X"33", X"36", X"33", X"1e", X"36", X"36", X"3c", X"23", X"0c", X"18", X"0c", X"00", X"7f", X"33", X"33", X"33", X"33", X"33", X"33", X"33", X"33", X"03", X"03", X"03", X"18", X"18", X"18", X"33", X"33", X"23", X"1b", X"1b", X"33", X"33", X"33", X"33", X"33", X"3c", X"33", X"33", X"33", X"03", X"36", X"36", X"1b", X"33", X"18", X"33", X"33", X"33", X"63", X"00", X"00", X"33", X"22", X"30", X"61", X"ce", X"1e", X"66", X"66", X"92", X"aa", X"6e", X"18", X"18", X"33", X"33", X"33", X"22", X"66", X"66", X"66", X"00", X"1e", X"0c", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"33", X"33", X"00", X"66", X"00", X"66", X"66", X"00", X"66", X"3e", X"63", X"36", X"23", X"23", X"23", X"00", X"0c", X"0c", X"0c", X"00", X"18", X"ff", X"ff", X"18", X"0c", X"00", X"33", X"1f", X"33", X"33", X"33", X"33", X"66", X"06", X"06", X"33", X"33", X"33", X"3c", X"0c", X"00", X"00", X"00", X"3f", X"1f", X"ce", X"e8", X"30", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"3f", X"00",
                                       X"00", X"7e", X"7e", X"08", X"00", X"7e", X"7e", X"00", X"00", X"00", X"00", X"1e", X"18", X"00", X"67", X"18", X"01", X"40", X"18", X"66", X"e8", X"63", X"7f", X"18", X"18", X"18", X"00", X"00", X"00", X"00", X"7f", X"08", X"00", X"0c", X"00", X"36", X"0c", X"31", X"6e", X"00", X"30", X"06", X"00", X"00", X"1c", X"00", X"1c", X"01", X"3e", X"3f", X"3f", X"1e", X"78", X"1e", X"1e", X"0c", X"1e", X"0e", X"00", X"18", X"30", X"00", X"06", X"0c", X"3e", X"33", X"3f", X"3c", X"1f", X"7f", X"0f", X"7c", X"33", X"1e", X"1e", X"67", X"7f", X"63", X"63", X"1c", X"0f", X"30", X"67", X"1e", X"1e", X"1e", X"0c", X"36", X"33", X"1e", X"7f", X"3c", X"40", X"3c", X"00", X"00", X"00", X"6e", X"3b", X"1e", X"6e", X"1e", X"0f", X"30", X"67", X"7e", X"33", X"67", X"7e", X"63", X"33", X"1e", X"3e", X"3e", X"0f", X"1e", X"1c", X"6e", X"0c", X"36", X"63", X"30", X"3f", X"38", X"18", X"07", X"00", X"00", X"1e", X"6e", X"1e", X"6e", X"6e", X"6e", X"6e", X"1e", X"3e", X"3e", X"3e", X"7e", X"7e", X"7e", X"33", X"33", X"3f", X"f7", X"7b", X"1e", X"1e", X"1e", X"6e", X"6e", X"30", X"1e", X"1e", X"1e", X"7f", X"1e", X"63", X"0e", X"6e", X"7e", X"1e", X"6e", X"33", X"63", X"00", X"00", X"1e", X"1c", X"00", X"30", X"fc", X"0c", X"cc", X"33", X"24", X"55", X"b6", X"18", X"18", X"33", X"33", X"33", X"1c", X"66", X"66", X"66", X"00", X"0c", X"0c", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"6e", X"33", X"00", X"66", X"00", X"66", X"66", X"00", X"66", X"63", X"3e", X"1f", X"3f", X"3f", X"3f", X"00", X"1e", X"1e", X"1e", X"00", X"18", X"ff", X"ff", X"18", X"1e", X"00", X"1e", X"03", X"1e", X"1e", X"1e", X"1e", X"ee", X"0f", X"0f", X"1e", X"1e", X"1e", X"30", X"1e", X"00", X"00", X"00", X"00", X"00", X"fc", X"e8", X"63", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                                       X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"00", X"00", X"00", X"00", X"00", X"00", X"7e", X"00", X"7e", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"78", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"ff", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"33", X"00", X"00", X"33", X"00", X"00", X"00", X"00", X"00", X"06", X"30", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"f8", X"c0", X"00", X"00", X"00", X"49", X"aa", X"eb", X"18", X"18", X"00", X"00", X"00", X"00", X"66", X"66", X"66", X"00", X"0c", X"00", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"00", X"00", X"00", X"66", X"00", X"66", X"66", X"00", X"66", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"ff", X"ff", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"18", X"00", X"00", X"00", X"00", X"00", X"00", X"c0", X"00", X"7e", X"00", X"0c", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
                                       X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"1e", X"00", X"00", X"1e", X"00", X"00", X"00", X"00", X"00", X"0f", X"78", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0f", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"06", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0f", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"92", X"55", X"6e", X"18", X"18", X"00", X"00", X"00", X"00", X"66", X"66", X"66", X"00", X"00", X"00", X"18", X"00", X"00", X"18", X"18", X"00", X"18", X"00", X"00", X"00", X"66", X"00", X"66", X"66", X"00", X"66", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"18", X"ff", X"ff", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"03", X"00", X"00", X"00", X"00", X"00", X"0f", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"0e", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00");


end fontROM;
