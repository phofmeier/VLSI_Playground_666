----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    17:42:44 01/08/2008
-- Design Name:
-- Module Name:    memory_int - Behavioral
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.std_logic_textio.all;
use std.textio.all;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memory_int is
   port ( clk  : in  std_logic;
          addr : in  std_logic_vector (10 downto 0);
          inp  : in  std_logic_vector (15 downto 0);
          outp : out std_logic_vector (15 downto 0);
          we   : in  std_logic);
end memory_int;


architecture Simulation of memory_int is
   type saveArray is array (0 to (2**addr'length-1)) of std_logic_vector(15 downto 0);
   signal data : saveArray := (others => (others => '0'));
begin

   mem_ctrl: process(clk)
      variable init : integer := 0;
      file inputfile : text open read_mode is "../memory.txt";
      variable inputline : line;
      variable inputval  : std_logic_vector(15 downto 0);
      variable address   : integer := 0;

   begin
      if init = 0 then
         while not endfile(inputfile) loop
            readline(inputfile, inputline);
            hread(inputline, inputval);
            data(address) <= inputval;
            address := address+1;
         end loop;
         init := 1;
      elsif rising_edge(clk) then
         if we = '1' then
            data(conv_integer(unsigned(addr))) <= inp;
            outp <= inp;
         else
            outp <= data(conv_integer(unsigned(addr)));
         end if;
      end if;
   end process mem_ctrl;
end Simulation;


architecture Synthesis of memory_int is
   type saveArray is array (0 to (2**addr'length-1)) of std_logic_vector(15 downto 0);
   signal data : saveArray := ( X"c008",
  X"c213",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"a200",
  X"8221",
  X"b000",
  X"8222",
  X"b005",
  X"8273",
  X"b001",
  X"821a",
  X"9265",
  X"8218",
  X"9262",
  X"9263",
  X"9264",
  X"9265",
  X"9266",
  X"9267",
  X"9268",
  X"9269",
  X"926a",
  X"926b",
  X"926c",
  X"f159",
  X"8262",
  X"d01d",
  X"f023",
  X"8218",
  X"9262",
  X"c01d",
  X"8265",
  X"d041",
  X"8262",
  X"2225",
  X"d04c",
  X"8262",
  X"2226",
  X"d04f",
  X"8262",
  X"2227",
  X"d058",
  X"8262",
  X"2234",
  X"d05b",
  X"8262",
  X"2229",
  X"d07e",
  X"8262",
  X"2235",
  X"d095",
  X"8265",
  X"2219",
  X"d04b",
  X"8262",
  X"222a",
  X"e04b",
  X"8233",
  X"2262",
  X"e04b",
  X"c084",
  X"8262",
  X"2228",
  X"d06b",
  X"8262",
  X"222a",
  X"e04b",
  X"8233",
  X"2262",
  X"e04b",
  X"c084",
  X"a100",
  X"8218",
  X"9263",
  X"c052",
  X"8219",
  X"9263",
  X"c052",
  X"8218",
  X"9265",
  X"f0cc",
  X"8263",
  X"9269",
  X"c0a7",
  X"8219",
  X"9264",
  X"c05d",
  X"821a",
  X"9264",
  X"8218",
  X"9265",
  X"826a",
  X"d064",
  X"f0c1",
  X"826f",
  X"c065",
  X"8266",
  X"9268",
  X"8218",
  X"9266",
  X"8264",
  X"926a",
  X"c0a7",
  X"8218",
  X"9265",
  X"8267",
  X"b021",
  X"8268",
  X"b021",
  X"8269",
  X"b021",
  X"826a",
  X"b021",
  X"8218",
  X"9267",
  X"9268",
  X"9269",
  X"926a",
  X"826b",
  X"1219",
  X"926b",
  X"c0a7",
  X"826b",
  X"d04b",
  X"8219",
  X"9265",
  X"f0e4",
  X"c0a7",
  X"821a",
  X"9265",
  X"8266",
  X"926d",
  X"821b",
  X"926e",
  X"f0f3",
  X"8262",
  X"222a",
  X"126f",
  X"9266",
  X"a004",
  X"3223",
  X"d0a7",
  X"8219",
  X"926c",
  X"c0a7",
  X"826b",
  X"d099",
  X"f0e4",
  X"c095",
  X"f0cc",
  X"8267",
  X"9266",
  X"826c",
  X"d09f",
  X"c0a7",
  X"f174",
  X"8246",
  X"b002",
  X"f1a5",
  X"f1c4",
  X"f174",
  X"f1b8",
  X"c0af",
  X"826c",
  X"d0bd",
  X"f174",
  X"8240",
  X"b002",
  X"f1a5",
  X"f174",
  X"f1b8",
  X"8218",
  X"9266",
  X"9267",
  X"9268",
  X"9269",
  X"926a",
  X"926b",
  X"926c",
  X"9265",
  X"821a",
  X"9265",
  X"8273",
  X"b001",
  X"a100",
  X"8262",
  X"9272",
  X"f183",
  X"a100",
  X"8266",
  X"926e",
  X"8268",
  X"926d",
  X"826a",
  X"2219",
  X"d0ca",
  X"f11f",
  X"c0cb",
  X"f0f3",
  X"a100",
  X"826a",
  X"d0d3",
  X"f0c1",
  X"826f",
  X"9266",
  X"8218",
  X"926a",
  X"8269",
  X"d0d9",
  X"8267",
  X"2266",
  X"9267",
  X"c0dc",
  X"8267",
  X"1266",
  X"9267",
  X"a004",
  X"3223",
  X"d0e1",
  X"8219",
  X"926c",
  X"8218",
  X"9266",
  X"a100",
  X"f0cc",
  X"8267",
  X"9266",
  X"a031",
  X"926a",
  X"a031",
  X"9269",
  X"a031",
  X"9268",
  X"a031",
  X"9267",
  X"826b",
  X"2219",
  X"926b",
  X"a100",
  X"8218",
  X"926f",
  X"9270",
  X"826d",
  X"e0f9",
  X"c0fe",
  X"5000",
  X"926d",
  X"8270",
  X"4000",
  X"9270",
  X"826e",
  X"e101",
  X"c106",
  X"5000",
  X"926e",
  X"8270",
  X"4000",
  X"9270",
  X"826e",
  X"d116",
  X"3219",
  X"d10e",
  X"826d",
  X"126f",
  X"e11c",
  X"926f",
  X"826d",
  X"126d",
  X"926d",
  X"e11c",
  X"826e",
  X"7000",
  X"926e",
  X"c107",
  X"8270",
  X"d11b",
  X"826f",
  X"5000",
  X"926f",
  X"a100",
  X"8219",
  X"926c",
  X"a100",
  X"8218",
  X"926f",
  X"9270",
  X"826d",
  X"e125",
  X"c12a",
  X"5000",
  X"926d",
  X"8270",
  X"4000",
  X"9270",
  X"826e",
  X"e12d",
  X"c132",
  X"5000",
  X"926e",
  X"8270",
  X"4000",
  X"9270",
  X"8219",
  X"9271",
  X"826d",
  X"226e",
  X"e13e",
  X"826e",
  X"126e",
  X"926e",
  X"8271",
  X"1271",
  X"9271",
  X"c134",
  X"826e",
  X"7000",
  X"926e",
  X"8271",
  X"7000",
  X"9271",
  X"d153",
  X"826d",
  X"226e",
  X"e14c",
  X"926d",
  X"8271",
  X"126f",
  X"926f",
  X"826e",
  X"7000",
  X"926e",
  X"8271",
  X"7000",
  X"9271",
  X"c144",
  X"8270",
  X"d158",
  X"826f",
  X"5000",
  X"926f",
  X"a100",
  X"f162",
  X"f1b8",
  X"825c",
  X"b002",
  X"f1a5",
  X"f174",
  X"f1b8",
  X"f174",
  X"a100",
  X"825d",
  X"b003",
  X"825e",
  X"9275",
  X"8237",
  X"b023",
  X"8275",
  X"2219",
  X"9275",
  X"d16d",
  X"c166",
  X"825d",
  X"9276",
  X"b003",
  X"8218",
  X"9278",
  X"9277",
  X"a100",
  X"8218",
  X"9277",
  X"9278",
  X"8276",
  X"125f",
  X"9276",
  X"b003",
  X"8260",
  X"2276",
  X"e17f",
  X"a100",
  X"825d",
  X"9276",
  X"b003",
  X"a100",
  X"8278",
  X"d19c",
  X"8272",
  X"121c",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"6000",
  X"9279",
  X"3239",
  X"b013",
  X"8219",
  X"9278",
  X"1277",
  X"9277",
  X"8261",
  X"2277",
  X"e19a",
  X"a100",
  X"f174",
  X"a100",
  X"8279",
  X"3272",
  X"b023",
  X"8218",
  X"9278",
  X"8219",
  X"1277",
  X"9277",
  X"a100",
  X"a012",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"7000",
  X"d1b7",
  X"9272",
  X"f183",
  X"a022",
  X"323b",
  X"d1b7",
  X"9272",
  X"f183",
  X"c1a5",
  X"a100",
  X"f174",
  X"825f",
  X"9275",
  X"8236",
  X"b023",
  X"8275",
  X"2219",
  X"9275",
  X"d1c2",
  X"c1bb",
  X"f174",
  X"a100",
  X"8218",
  X"927a",
  X"927b",
  X"927c",
  X"927d",
  X"927e",
  X"8266",
  X"e20c",
  X"8266",
  X"221d",
  X"9266",
  X"e1d4",
  X"827a",
  X"1219",
  X"927a",
  X"c1cc",
  X"121d",
  X"221e",
  X"9266",
  X"e1dd",
  X"827b",
  X"1219",
  X"927b",
  X"8266",
  X"c1d5",
  X"121e",
  X"221f",
  X"9266",
  X"e1e6",
  X"827c",
  X"1219",
  X"927c",
  X"8266",
  X"c1de",
  X"121f",
  X"2220",
  X"9266",
  X"e1ef",
  X"827d",
  X"1219",
  X"927d",
  X"8266",
  X"c1e7",
  X"1220",
  X"927e",
  X"827a",
  X"d1fd",
  X"f208",
  X"827b",
  X"f208",
  X"827c",
  X"f208",
  X"827d",
  X"f208",
  X"827b",
  X"f208",
  X"a100",
  X"827b",
  X"d200",
  X"c1f5",
  X"827c",
  X"d203",
  X"c1f7",
  X"827d",
  X"d206",
  X"c1f9",
  X"827e",
  X"c1fb",
  X"1238",
  X"9272",
  X"f183",
  X"a100",
  X"5000",
  X"9266",
  X"8226",
  X"9272",
  X"f183",
  X"8266",
  X"c1cc",
  X"b030",
  X"8fff",
  X"9262",
  X"a020",
  X"a200",
  X"0000",
  X"0001",
  X"0002",
  X"000a",
  X"ff00",
  X"2710",
  X"03e8",
  X"0064",
  X"000a",
  X"07ff",
  X"0102",
  X"0008",
  X"00ff",
  X"002b",
  X"002d",
  X"002a",
  X"0028",
  X"0029",
  X"0030",
  X"0031",
  X"0032",
  X"0033",
  X"0034",
  X"0035",
  X"0036",
  X"0037",
  X"0038",
  X"0039",
  X"002f",
  X"003d",
  X"2d2d",
  X"2020",
  X"0030",
  X"ff20",
  X"ff00",
  X"00ff",
  X"4572",
  X"726f",
  X"7221",
  X"0000",
  X"023c",
  X"5265",
  X"7375",
  X"6c74",
  X"3a20",
  X"0000",
  X"0241",
  X"5765",
  X"6c63",
  X"6f6d",
  X"6520",
  X"746f",
  X"2074",
  X"6865",
  X"2075",
  X"6c74",
  X"696d",
  X"6174",
  X"6520",
  X"4c4d",
  X"4520",
  X"6361",
  X"6c63",
  X"756c",
  X"6174",
  X"6f72",
  X"2120",
  X"0000",
  X"0247",
  X"0800",
  X"0640",
  X"0028",
  X"0e40",
  X"004f",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0274",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  X"0000",
  others => X"0000" );
begin

   mem_ctrl: process(clk)
   begin
      if rising_edge(clk) then
         if we = '1' then
            data(conv_integer(unsigned(addr))) <= inp;
            outp <= inp;
         else
            outp <= data(conv_integer(unsigned(addr)));
         end if;
      end if;
   end process mem_ctrl;
end Synthesis;







